library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.NUMERIC_STD.all;

entity RotateRightOp is
Port (A : in std_logic_vector(15 downto 0);
rorEn: in std_logic;
Result : out std_logic_vector(15 downto 0));
end RotateRightOp;

architecture Behavioral of RotateRightOp is

signal Output: std_logic_vector(15 downto 0);

begin

Output <= std_logic_vector(unsigned(A) ror 1);

process(Output, rorEn)
begin

if rorEn ='1' then
   Result <= Output;
else Result <= "ZZZZZZZZZZZZZZZZ";
end if;
end process;

end Behavioral;
